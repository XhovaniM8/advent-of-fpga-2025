module counter (
    input logic clk,
    input logic rst,
    output logic [7:0] count
);
    always_ff @(posedge clk or posedge rst)
        if (rst) count <= 8'h0;
        else count <= count + 1'b1;
endmodule
